module Fetch (
    
);
endmodule